module SubWord(
	input wire [7:0] S0_in,
	input wire [7:0] S1_in,
	input wire [7:0] S2_in,
	input wire [7:0] S3_in,
	output wire [7:0] D0_out,
	output wire [7:0] D1_out,
	output wire [7:0] D2_out,
	output wire [7:0] D3_out	
	);
	
	sbox sb0 (.S_in(S0_in), .D_out(D0_out));
	sbox sb1 (.S_in(S1_in), .D_out(D1_out));
	sbox sb2 (.S_in(S2_in), .D_out(D2_out));
	sbox sb3 (.S_in(S3_in), .D_out(D3_out));
	
endmodule

module sbox(
	input  wire   [7:0] S_in,
    output reg    [7:0] D_out);
                  
always @*
begin
    case (S_in)
       8'h00: D_out = 8'h63;
	   8'h01: D_out = 8'h7c;
	   8'h02: D_out = 8'h77;
	   8'h03: D_out = 8'h7b;
	   8'h04: D_out = 8'hf2;
	   8'h05: D_out = 8'h6b;
	   8'h06: D_out = 8'h6f;
	   8'h07: D_out = 8'hc5;
	   8'h08: D_out = 8'h30;
	   8'h09: D_out = 8'h01;
	   8'h0a: D_out = 8'h67;
	   8'h0b: D_out = 8'h2b;
	   8'h0c: D_out = 8'hfe;
	   8'h0d: D_out = 8'hd7;
	   8'h0e: D_out = 8'hab;
	   8'h0f: D_out = 8'h76;
	   8'h10: D_out = 8'hca;
	   8'h11: D_out = 8'h82;
	   8'h12: D_out = 8'hc9;
	   8'h13: D_out = 8'h7d;
	   8'h14: D_out = 8'hfa;
	   8'h15: D_out = 8'h59;
	   8'h16: D_out = 8'h47;
	   8'h17: D_out = 8'hf0;
	   8'h18: D_out = 8'had;
	   8'h19: D_out = 8'hd4;
	   8'h1a: D_out = 8'ha2;
	   8'h1b: D_out = 8'haf;
	   8'h1c: D_out = 8'h9c;
	   8'h1d: D_out = 8'ha4;
	   8'h1e: D_out = 8'h72;
	   8'h1f: D_out = 8'hc0;
	   8'h20: D_out = 8'hb7;
	   8'h21: D_out = 8'hfd;
	   8'h22: D_out = 8'h93;
	   8'h23: D_out = 8'h26;
	   8'h24: D_out = 8'h36;
	   8'h25: D_out = 8'h3f;
	   8'h26: D_out = 8'hf7;
	   8'h27: D_out = 8'hcc;
	   8'h28: D_out = 8'h34;
	   8'h29: D_out = 8'ha5;
	   8'h2a: D_out = 8'he5;
	   8'h2b: D_out = 8'hf1;
	   8'h2c: D_out = 8'h71;
	   8'h2d: D_out = 8'hd8;
	   8'h2e: D_out = 8'h31;
	   8'h2f: D_out = 8'h15;
	   8'h30: D_out = 8'h04;
	   8'h31: D_out = 8'hc7;
	   8'h32: D_out = 8'h23;
	   8'h33: D_out = 8'hc3;
	   8'h34: D_out = 8'h18;
	   8'h35: D_out = 8'h96;
	   8'h36: D_out = 8'h05;
	   8'h37: D_out = 8'h9a;
	   8'h38: D_out = 8'h07;
	   8'h39: D_out = 8'h12;
	   8'h3a: D_out = 8'h80;
	   8'h3b: D_out = 8'he2;
	   8'h3c: D_out = 8'heb;
	   8'h3d: D_out = 8'h27;
	   8'h3e: D_out = 8'hb2;
	   8'h3f: D_out = 8'h75;
	   8'h40: D_out = 8'h09;
	   8'h41: D_out = 8'h83;
	   8'h42: D_out = 8'h2c;
	   8'h43: D_out = 8'h1a;
	   8'h44: D_out = 8'h1b;
	   8'h45: D_out = 8'h6e;
	   8'h46: D_out = 8'h5a;
	   8'h47: D_out = 8'ha0;
	   8'h48: D_out = 8'h52;
	   8'h49: D_out = 8'h3b;
	   8'h4a: D_out = 8'hd6;
	   8'h4b: D_out = 8'hb3;
	   8'h4c: D_out = 8'h29;
	   8'h4d: D_out = 8'he3;
	   8'h4e: D_out = 8'h2f;
	   8'h4f: D_out = 8'h84;
	   8'h50: D_out = 8'h53;
	   8'h51: D_out = 8'hd1;
	   8'h52: D_out = 8'h00;
	   8'h53: D_out = 8'hed;
	   8'h54: D_out = 8'h20;
	   8'h55: D_out = 8'hfc;
	   8'h56: D_out = 8'hb1;
	   8'h57: D_out = 8'h5b;
	   8'h58: D_out = 8'h6a;
	   8'h59: D_out = 8'hcb;
	   8'h5a: D_out = 8'hbe;
	   8'h5b: D_out = 8'h39;
	   8'h5c: D_out = 8'h4a;
	   8'h5d: D_out = 8'h4c;
	   8'h5e: D_out = 8'h58;
	   8'h5f: D_out = 8'hcf;
	   8'h60: D_out = 8'hd0;
	   8'h61: D_out = 8'hef;
	   8'h62: D_out = 8'haa;
	   8'h63: D_out = 8'hfb;
	   8'h64: D_out = 8'h43;
	   8'h65: D_out = 8'h4d;
	   8'h66: D_out = 8'h33;
	   8'h67: D_out = 8'h85;
	   8'h68: D_out = 8'h45;
	   8'h69: D_out = 8'hf9;
	   8'h6a: D_out = 8'h02;
	   8'h6b: D_out = 8'h7f;
	   8'h6c: D_out = 8'h50;
	   8'h6d: D_out = 8'h3c;
	   8'h6e: D_out = 8'h9f;
	   8'h6f: D_out = 8'ha8;
	   8'h70: D_out = 8'h51;
	   8'h71: D_out = 8'ha3;
	   8'h72: D_out = 8'h40;
	   8'h73: D_out = 8'h8f;
	   8'h74: D_out = 8'h92;
	   8'h75: D_out = 8'h9d;
	   8'h76: D_out = 8'h38;
	   8'h77: D_out = 8'hf5;
	   8'h78: D_out = 8'hbc;
	   8'h79: D_out = 8'hb6;
	   8'h7a: D_out = 8'hda;
	   8'h7b: D_out = 8'h21;
	   8'h7c: D_out = 8'h10;
	   8'h7d: D_out = 8'hff;
	   8'h7e: D_out = 8'hf3;
	   8'h7f: D_out = 8'hd2;
	   8'h80: D_out = 8'hcd;
	   8'h81: D_out = 8'h0c;
	   8'h82: D_out = 8'h13;
	   8'h83: D_out = 8'hec;
	   8'h84: D_out = 8'h5f;
	   8'h85: D_out = 8'h97;
	   8'h86: D_out = 8'h44;
	   8'h87: D_out = 8'h17;
	   8'h88: D_out = 8'hc4;
	   8'h89: D_out = 8'ha7;
	   8'h8a: D_out = 8'h7e;
	   8'h8b: D_out = 8'h3d;
	   8'h8c: D_out = 8'h64;
	   8'h8d: D_out = 8'h5d;
	   8'h8e: D_out = 8'h19;
	   8'h8f: D_out = 8'h73;
	   8'h90: D_out = 8'h60;
	   8'h91: D_out = 8'h81;
	   8'h92: D_out = 8'h4f;
	   8'h93: D_out = 8'hdc;
	   8'h94: D_out = 8'h22;
	   8'h95: D_out = 8'h2a;
	   8'h96: D_out = 8'h90;
	   8'h97: D_out = 8'h88;
	   8'h98: D_out = 8'h46;
	   8'h99: D_out = 8'hee;
	   8'h9a: D_out = 8'hb8;
	   8'h9b: D_out = 8'h14;
	   8'h9c: D_out = 8'hde;
	   8'h9d: D_out = 8'h5e;
	   8'h9e: D_out = 8'h0b;
	   8'h9f: D_out = 8'hdb;
	   8'ha0: D_out = 8'he0;
	   8'ha1: D_out = 8'h32;
	   8'ha2: D_out = 8'h3a;
	   8'ha3: D_out = 8'h0a;
	   8'ha4: D_out = 8'h49;
	   8'ha5: D_out = 8'h06;
	   8'ha6: D_out = 8'h24;
	   8'ha7: D_out = 8'h5c;
	   8'ha8: D_out = 8'hc2;
	   8'ha9: D_out = 8'hd3;
	   8'haa: D_out = 8'hac;
	   8'hab: D_out = 8'h62;
	   8'hac: D_out = 8'h91;
	   8'had: D_out = 8'h95;
	   8'hae: D_out = 8'he4;
	   8'haf: D_out = 8'h79;
	   8'hb0: D_out = 8'he7;
	   8'hb1: D_out = 8'hc8;
	   8'hb2: D_out = 8'h37;
	   8'hb3: D_out = 8'h6d;
	   8'hb4: D_out = 8'h8d;
	   8'hb5: D_out = 8'hd5;
	   8'hb6: D_out = 8'h4e;
	   8'hb7: D_out = 8'ha9;
	   8'hb8: D_out = 8'h6c;
	   8'hb9: D_out = 8'h56;
	   8'hba: D_out = 8'hf4;
	   8'hbb: D_out = 8'hea;
	   8'hbc: D_out = 8'h65;
	   8'hbd: D_out = 8'h7a;
	   8'hbe: D_out = 8'hae;
	   8'hbf: D_out = 8'h08;
	   8'hc0: D_out = 8'hba;
	   8'hc1: D_out = 8'h78;
	   8'hc2: D_out = 8'h25;
	   8'hc3: D_out = 8'h2e;
	   8'hc4: D_out = 8'h1c;
	   8'hc5: D_out = 8'ha6;
	   8'hc6: D_out = 8'hb4;
	   8'hc7: D_out = 8'hc6;
	   8'hc8: D_out = 8'he8;
	   8'hc9: D_out = 8'hdd;
	   8'hca: D_out = 8'h74;
	   8'hcb: D_out = 8'h1f;
	   8'hcc: D_out = 8'h4b;
	   8'hcd: D_out = 8'hbd;
	   8'hce: D_out = 8'h8b;
	   8'hcf: D_out = 8'h8a;
	   8'hd0: D_out = 8'h70;
	   8'hd1: D_out = 8'h3e;
	   8'hd2: D_out = 8'hb5;
	   8'hd3: D_out = 8'h66;
	   8'hd4: D_out = 8'h48;
	   8'hd5: D_out = 8'h03;
	   8'hd6: D_out = 8'hf6;
	   8'hd7: D_out = 8'h0e;
	   8'hd8: D_out = 8'h61;
	   8'hd9: D_out = 8'h35;
	   8'hda: D_out = 8'h57;
	   8'hdb: D_out = 8'hb9;
	   8'hdc: D_out = 8'h86;
	   8'hdd: D_out = 8'hc1;
	   8'hde: D_out = 8'h1d;
	   8'hdf: D_out = 8'h9e;
	   8'he0: D_out = 8'he1;
	   8'he1: D_out = 8'hf8;
	   8'he2: D_out = 8'h98;
	   8'he3: D_out = 8'h11;
	   8'he4: D_out = 8'h69;
	   8'he5: D_out = 8'hd9;
	   8'he6: D_out = 8'h8e;
	   8'he7: D_out = 8'h94;
	   8'he8: D_out = 8'h9b;
	   8'he9: D_out = 8'h1e;
	   8'hea: D_out = 8'h87;
	   8'heb: D_out = 8'he9;
	   8'hec: D_out = 8'hce;
	   8'hed: D_out = 8'h55;
	   8'hee: D_out = 8'h28;
	   8'hef: D_out = 8'hdf;
	   8'hf0: D_out = 8'h8c;
	   8'hf1: D_out = 8'ha1;
	   8'hf2: D_out = 8'h89;
	   8'hf3: D_out = 8'h0d;
	   8'hf4: D_out = 8'hbf;
	   8'hf5: D_out = 8'he6;
	   8'hf6: D_out = 8'h42;
	   8'hf7: D_out = 8'h68;
	   8'hf8: D_out = 8'h41;
	   8'hf9: D_out = 8'h99;
	   8'hfa: D_out = 8'h2d;
	   8'hfb: D_out = 8'h0f;
	   8'hfc: D_out = 8'hb0;
	   8'hfd: D_out = 8'h54;
	   8'hfe: D_out = 8'hbb;
	   8'hff: D_out = 8'h16;
	endcase
end
endmodule
